library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity display_seven_seg is
    Port ( clock_in : in STD_LOGIC; -- 100 MHz input clock
           reset_timer : in STD_LOGIC; -- Reset signal (Resetting the internal signals to known states)
           d0: in std_logic_vector(3 downto 0);
           d1: in std_logic_vector(3 downto 0);
           d2: in std_logic_vector(3 downto 0);
           d3: in std_logic_vector(3 downto 0);
           an : out STD_LOGIC_VECTOR (3 downto 0); -- Anodes signal for display
           seg : out STD_LOGIC_VECTOR (6 downto 0) -- Cathodes signal for display
           );
end display_seven_seg;

architecture Behavioral of display_seven_seg is
    
    component Timing_block is
        Port (
            clk_in : in STD_LOGIC; -- 100 MHz input clock
            reset : in STD_LOGIC; -- Reset signal (Resetting the internal signals to known states)
            mux_select : out STD_LOGIC_VECTOR (1 downto 0); -- Signal for the mux
            anodes_tout : out STD_LOGIC_VECTOR (3 downto 0); -- Anodes signal for display
        );
    end component;

    component seven_seg_decoder_decimal is
        port (
            dec_in : in std_logic_vector(3 downto 0);
            dec_out : out std_logic_vector(6 downto 0)
        );
    end component;

    component MUX_4BIT is
        port(
            mux_s : in std_logic_vector(1 downto 0);
            mux_d0 : in std_logic_vector(3 downto 0);
            mux_d1 : in std_logic_vector(3 downto 0);
            mux_d2 : in std_logic_vector(3 downto 0);
            mux_d3 : in std_logic_vector(3 downto 0);
            mux_out_to : out std_logic_vector(3 downto 0);
        );
    end component;
    
    signal mux_sel: std_logic_vector(1 downto 0);
    signal mux_out_dec: std_logic_vector(3 downto 0);
    
begin
    Timer_Block : Timing_Block port map (clock_in,reset_timer,mux_sel,an);
    MUX_Block : MUX_4BIT port map (mux_sel,d0,d1,d2,d3,mux_out_dec);
    Decoder_Block : seven_seg_decoder_decimal port map (mux_out_dec,seg);  

end Behavioral;
